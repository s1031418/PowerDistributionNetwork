# R=RESISTANCE RPERSQ* L/W
RVDD3_1 M5_0_1000000  M5_277600_1000000 1.1104
RVDD3_2 M5_277600_1000000  M6_277600_1000000 1.0
RVDD3_3 M6_277600_1000000  M6_277600_1896600  1.8032
RVDD3_4 M6_277600_1896600 M6_1543000_1896600  2.5508
RVDD3_5 M5_277600_1000000 M5_277600_316600    2.7736
RVDD3_6 M5_277600_316600  M5_391000_316600   0.4936
V_VDD3_1 M5_0_1000000 gnd 1.0
I_VDD3_1 M6_1543000_1896600 gnd  3e-3
I_VDD3_2 M5_391000_316600   gnd 2e-3

RVDD2_1 M5_0_500000 M5_113700_500000   0.4548
RVDD2_2 M5_113700_500000 M6_113700_500000   1.0
RVDD2_3 M6_113700_500000 M6_113700_547900  0.1058
RVDD2_4 M6_113700_547900 M6_1701000_547900  3.1946
V_VDD2_1 M5_0_500000 gnd 1.0
I_VDD2_1 M6_1701000_547900 gnd 2e-3

RVDD1_1 M6_200000_0 M6_200000_180600  0.3612
RVDD1_2 M6_200000_180600 M6_1611500_180600   2.833
RVDD1_3 M6_1611500_180600 M6_1611500_367500  0.3938
RVDD1_4 M6_1611500_367500 M6_1701000_367500  0.199
V_VDD1_1 M6_200000_0 gnd 1.0
I_VDD1_1 M6_1701000_367500 gnd 5e-3

.tran 1ns 1ns
.end
