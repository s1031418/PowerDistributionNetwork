#Comments
RVDD1_1 METAL6_200000_175600 METAL6_1606500_175600 1.4065
RVDD1_2 METAL6_200000_0 METAL6_200000_175600 0.1756
RVDD1_3 METAL6_1606500_362500 METAL6_1701000_379000 0.0945
RVDD1_4 METAL6_1606500_175600 METAL6_1606500_362500 0.1869
V_VDD1_1 METAL6_200000_0 gnd 1.0
IVDD1_1 METAL6_1701000_379000 gnd 0.005000

RVDD2_1 METAL5_0_500000 METAL5_108700_500000 0.4348
RVDD2_2 METAL6_108700_542900 METAL6_1701000_569000 3.1846
RVDD2_3 METAL6_108700_500000 METAL6_108700_542900 0.0858
RVDD2_4 METAL5_108700_500000 METAL6_108700_500000 1
V_VDD2_1 METAL5_0_500000 gnd 1.0
IVDD2_1 METAL6_1701000_569000 gnd 0.002000

RVDD3_1 METAL5_0_1000000 METAL5_272600_1000000 1.0904
RVDD3_2 METAL5_272600_316600 METAL5_391000_345000 0.4736
RVDD3_3 METAL6_272600_1879600 METAL6_1543000_1919000 2.5408
RVDD3_4 METAL6_272600_1891600 METAL6_1543000_1919000 2.5408
RVDD3_5 METAL6_272600_1903600 METAL6_1543000_1919000 2.5408
RVDD3_6 METAL5_272600_316600 METAL5_272600_1000000 2.7336
RVDD3_7 METAL6_272600_1000000 METAL6_272600_1879600 1.7592
RVDD3_8 METAL6_272600_1879600 METAL6_272600_1891600 0.024
RVDD3_9 METAL6_272600_1891600 METAL6_272600_1903600 0.024
RVDD3_10 METAL5_272600_1000000 METAL6_272600_1000000 1
V_VDD3_1 METAL5_0_1000000 gnd 1.0
IVDD3_1 METAL5_391000_345000 gnd 0.002000
IVDD3_2 METAL6_1543000_1919000 gnd 0.003000

.tran 1ns 1ns
.end
.control
set noaskquit
run
quit
.enddc
