module top (VDD1, VDD2, VDD3, VDD4, VDD5, VDD6, VDD7, VDD8, VDD9, VDD10, VDD11, VDD12, VDD13, VDD14, VDD15, VDD16, VDD17, VDD18, VDD19, VDD20, VDD21, VDD22, VDD23, VDD24, VDD25, VDD26, VDD_111a, VDD_111b );
  input VDD1, VDD2, VDD3, VDD4, VDD5, VDD6, VDD7, VDD8, VDD9, VDD10, VDD11, VDD12, VDD13, VDD14, VDD15, VDD16, VDD17, VDD18, VDD19, VDD20, VDD21, VDD22, VDD23, VDD24, VDD25, VDD26, VDD_111a, VDD_111b ;


/* multi-in-a */
  block6 B6_01 ( .VDD_A(VDD_111a) );
  block6 B6_02 ( .VDD_A(VDD_111a) );
  block6 B6_03 ( .VDD_A(VDD_111a) );

// multi-in-b
  block6 B6_04 ( .VDD_A(VDD_111b) );
  block6 B6_05 ( .VDD_A(VDD_111b) );
  block6 B6_06 ( .VDD_A(VDD_111b) );
 



endmodule

