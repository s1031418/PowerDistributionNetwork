
module top (VDD1, VDD2, VDD3, VDD4, VDD5);
  input VDD1, VDD2, VDD3, VDD4, VDD5;

  block9 B_T0 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5) );
  block9 B_T1 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_T2 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_T3 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_T4 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_T5 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_T6 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_T7 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_T8 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_T9 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_B0 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_B1 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_B2 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_B3 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_B4 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_B5 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_B6 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_B7 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_B8 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
  block9 B_B9 ( .VDD_A(VDD1), .VDD_B(VDD2), .VDD_C(VDD3), .VDD_D(VDD4), .VDD_E(VDD5)  );
endmodule

