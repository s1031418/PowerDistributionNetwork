# R=RESISTANCE RPERSQ* L/W
RVDD1_1 M6_200000_0 M6_200000_185600  0.1856
RVDD1_2 M6_200000_185600 M6_1616500_175600   1.4265
RVDD1_3 M6_1616500_175600 M6_1606500_372500  0.2069
RVDD1_4 M6_1606500_372500 M6_1701000_362500  0.1045
V_VDD1_1 M6_200000_0 gnd 1.0
I_VDD1_1 M6_1701000_362500 gnd 5e-3

RVDD2_1 M5_0_500000 M5_113700_500000 0.4548
RVDD2_2 M5_113700_500000 M6_108700_500000 1.0
RVDD2_3 M6_108700_500000 M6_108700_547900 0.1058
RVDD2_4 M6_108700_547900 M6_1701000_542900 3.1946
V_VDD2_1 M5_0_500000 gnd 1.0
I_VDD2_1 M6_1701000_542900 gnd 2e-3

RVDD3_1 M5_0_1000000  M5_277600_1000000 1.1104
RVDD3_2 M5_277600_1000000 M5_272600_316600 2.7736
RVDD3_3 M5_272600_316600  M5_391000_316600 0.4936
RVDD3_4 M5_277600_1000000  M6_272600_1000000 1.0
RVDD3_5 M6_272600_1000000 M6_272600_1884600 1.7792
RVDD3_6 M6_272600_1884600 M6_272600_1896600 0.024
RVDD3_7 M6_272600_1896600 M6_272600_1908600 0.024
RVDD3_8 M6_272600_1884600  M6_1543000_1879600 2.5508
RVDD3_9 M6_272600_1896600  M6_1543000_1879600 2.5508
RVDD3_10 M6_272600_1908600  M6_1543000_1879600 2.5508
V_VDD3_1 M5_0_1000000 gnd 1.0
I_VDD3_1 M6_1543000_1879600  gnd  3e-3
I_VDD3_2 M5_391000_316600   gnd 2e-3

.tran 1ns 1ns
.end
