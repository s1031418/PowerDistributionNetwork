VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
#BUSBITCHARS "d" ;
#DIVIDERCHAR "/" ;

SITE unit
  CLASS CORE ;
  SYMMETRY X Y ;
  SIZE 0.2 BY 1.8 ;
END unit


MACRO block1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 800 BY 500 ;
  SYMMETRY X Y R90 ;

  PIN VDD_A
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    LAYER METAL5 ;
       RECT 0 10 5 60 ;
    LAYER METAL6 ;
       RECT 0 10 5 60 ;
    END 
  END VDD_A
  PIN VDD_B
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    LAYER METAL5 ;
       RECT 0 200 5 250 ;
    LAYER METAL6 ;
       RECT 0 200 5 250 ;
    END
  END VDD_B

  OBS
    LAYER METAL1 ;
       RECT 0 0 800 500 ;
    LAYER METAL2 ;
       RECT 0 0 800 500 ;
    LAYER METAL3 ;
       RECT 0 0 800 500 ;
    LAYER METAL4 ;
       RECT 0 0 800 500 ;
    LAYER METAL5 ;
       RECT 0 0 800 500 ;
    LAYER METAL6 ;
       RECT 0 0 800 500 ;
  END
END block1

MACRO block2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 50 BY 300 ;
  SYMMETRY X Y R90 ;

  PIN VDD_A
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    LAYER METAL5 ;
       RECT 0 50 5 70 ;
    LAYER METAL6 ;
       RECT 0 50 5 70 ;
    END
  END VDD_A

  OBS
    LAYER METAL1 ;
       RECT 0 0 50 300 ;
    LAYER METAL2 ;
       RECT 0 0 50 300 ;
    LAYER METAL3 ;
       RECT 0 0 50 300 ;
    LAYER METAL4 ;
       RECT 0 0 50 300 ;
    LAYER METAL5 ;
       RECT 0 0 50 300 ;
    LAYER METAL6 ;
       RECT 0 0 50 300 ;
  END  
END block2

MACRO block3
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 100 BY 200 ;
  SYMMETRY X Y R90 ;

  PIN VDD_A
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    LAYER METAL2 ;
       RECT 0 50 5 70 ;
    LAYER METAL3 ;
       RECT 0 50 5 70 ;
    END
  END VDD_A

  OBS
    LAYER METAL1 ;
       RECT 0 0 100 200 ;
    LAYER METAL2 ;
       RECT 0 0 100 200 ;
    LAYER METAL3 ;
       RECT 0 0 100 200 ;
  END
END block3

MACRO block4
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 300 BY 300 ;
  SYMMETRY X Y R90 ;

  PIN VDD_A
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    LAYER METAL5 ;
       RECT 0 100 5 200 ;
    LAYER METAL6 ;
       RECT 0 100 5 200 ;
    END
  END VDD_A

  OBS
    LAYER METAL1 ;
       RECT 0 0 300 300 ;
    LAYER METAL2 ;
       RECT 0 0 300 300 ;
    LAYER METAL3 ;
       RECT 0 0 300 300 ;
    LAYER METAL4 ;
       RECT 0 0 300 300 ;
    LAYER METAL5 ;
       RECT 0 0 300 300 ;
    LAYER METAL6 ;
       RECT 0 0 300 300 ;
  END
END block4

MACRO block5
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 250 BY 700 ;
  SYMMETRY X Y R90 ;

  PIN VDD_A
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    LAYER METAL5 ;
       RECT 0 150 5 180 ;
    LAYER METAL6 ;
       RECT 0 150 5 180 ;
    END
  END VDD_A
  PIN VDD_B
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    LAYER METAL5 ;
       RECT 0 250 5 280 ;
    LAYER METAL6 ;
       RECT 0 250 5 280 ;
    END
  END VDD_B
  PIN VDD_C
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    LAYER METAL5 ;
       RECT 0 350 5 380 ;
    LAYER METAL6 ;
       RECT 0 350 5 380 ;
    END
  END VDD_C
  PIN VDD_D
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    LAYER METAL5 ;
       RECT 0 450 5 480 ;
    LAYER METAL6 ;
       RECT 0 450 5 480 ;
    END
  END VDD_D
  PIN VDD_E
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    LAYER METAL5 ;
       RECT 0 550 5 580 ;
    LAYER METAL6 ;
       RECT 0 550 5 580 ;
    END
  END VDD_E

  OBS
    LAYER METAL1 ;
       RECT 0 0 250 700 ;
    LAYER METAL2 ; 
       RECT 0 0 250 700 ;
    LAYER METAL3 ; 
       RECT 0 0 250 700 ;
    LAYER METAL4 ;
       RECT 0 0 250 700 ;
    LAYER METAL5 ;
       RECT 0 0 250 700 ;
    LAYER METAL6 ;
       RECT 0 0 250 700 ;
  END  
END block5

END LIBRARY
